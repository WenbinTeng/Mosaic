`timescale 1ns/1ps

module top (
    input clk_100MHz,
    input aresetn
);
    
endmodule